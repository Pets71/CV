--Package for defining the enum operation to all.
package operation_package is
    type op_type is 
        (ADD, COM, DEC, INC, SUB, BSF, BCF, ANP, IOR, XOP, SWP, RLF, RRF, MOV, CLR, NOP);
end operation_package;



